// Compiler Directives

// Used for extra debug outputs for the LED display, turn on for FPGA prototyping, off for simulation
`define VALIDATION 1