module partial_product (
  input  [31:0] a, b,  
  output [31:0] pp0,  pp1,  pp2,  pp3,  pp4,  pp5,  pp6,  pp7, 
                pp8,  pp9,  pp10, pp11, pp12, pp13, pp14, pp15,
                pp16, pp17, pp18, pp19, pp20, pp21, pp22, pp23, 
                pp24, pp25, pp26, pp27, pp28, pp29, pp30, pp31);

/*
 Better way w/ looping
( input  logic [31:0] A, B;
  output logic [31:0] PP [31:0] ); 
  
  always_comb begin
    // For each PP
    for (int index=0; index<32; index++) begin
      // For each bit of PP
      for (int a_bit=0; a_bit<32; a_bit++) begin
        // For each bit of B
        for (int b_bit=0; b_bit<32; b_bit++) begin
          // AND current bit of A with bit of B corresponding to index of PP
          PP[index][a_bit] = A[a_bit] & B[b_bit];
        end
      end
    end
  end
*/
  
    assign pp0[0]   = a[0]  & b[0];
    assign pp1[0]   = a[0]  & b[1];
    assign pp2[0]   = a[0]  & b[2];
    assign pp3[0]   = a[0]  & b[3];
    assign pp4[0]   = a[0]  & b[4];
    assign pp5[0]   = a[0]  & b[5];
    assign pp6[0]   = a[0]  & b[6];
    assign pp7[0]   = a[0]  & b[7];
    assign pp8[0]   = a[0]  & b[8];
    assign pp9[0]   = a[0]  & b[9];
    assign pp10[0]  = a[0]  & b[10];
    assign pp11[0]  = a[0]  & b[11];
    assign pp12[0]  = a[0]  & b[12];
    assign pp13[0]  = a[0]  & b[13];
    assign pp14[0]  = a[0]  & b[14];
    assign pp15[0]  = a[0]  & b[15];
    assign pp16[0]  = a[0]  & b[16];
    assign pp17[0]  = a[0]  & b[17];
    assign pp18[0]  = a[0]  & b[18];
    assign pp19[0]  = a[0]  & b[19];
    assign pp20[0]  = a[0]  & b[20];
    assign pp21[0]  = a[0]  & b[21];
    assign pp22[0]  = a[0]  & b[22];
    assign pp23[0]  = a[0]  & b[23];
    assign pp24[0]  = a[0]  & b[24];
    assign pp25[0]  = a[0]  & b[25];
    assign pp26[0]  = a[0]  & b[26];
    assign pp27[0]  = a[0]  & b[27];
    assign pp28[0]  = a[0]  & b[28];
    assign pp29[0]  = a[0]  & b[29];
    assign pp30[0]  = a[0]  & b[30];
    assign pp31[0]  = a[0]  & b[31];

    assign pp0[1]   = a[1]  & b[0];
    assign pp1[1]   = a[1]  & b[1];
    assign pp2[1]   = a[1]  & b[2];
    assign pp3[1]   = a[1]  & b[3];
    assign pp4[1]   = a[1]  & b[4];
    assign pp5[1]   = a[1]  & b[5];
    assign pp6[1]   = a[1]  & b[6];
    assign pp7[1]   = a[1]  & b[7];
    assign pp8[1]   = a[1]  & b[8];
    assign pp9[1]   = a[1]  & b[9];
    assign pp10[1]  = a[1]  & b[10];
    assign pp11[1]  = a[1]  & b[11];
    assign pp12[1]  = a[1]  & b[12];
    assign pp13[1]  = a[1]  & b[13];
    assign pp14[1]  = a[1]  & b[14];
    assign pp15[1]  = a[1]  & b[15];
    assign pp16[1]  = a[1]  & b[16];
    assign pp17[1]  = a[1]  & b[17];
    assign pp18[1]  = a[1]  & b[18];
    assign pp19[1]  = a[1]  & b[19];
    assign pp20[1]  = a[1]  & b[20];
    assign pp21[1]  = a[1]  & b[21];
    assign pp22[1]  = a[1]  & b[22];
    assign pp23[1]  = a[1]  & b[23];
    assign pp24[1]  = a[1]  & b[24];
    assign pp25[1]  = a[1]  & b[25];
    assign pp26[1]  = a[1]  & b[26];
    assign pp27[1]  = a[1]  & b[27];
    assign pp28[1]  = a[1]  & b[28];
    assign pp29[1]  = a[1]  & b[29];
    assign pp30[1]  = a[1]  & b[30];
    assign pp31[1]  = a[1]  & b[31];

    assign pp0[2]   = a[2]  & b[0];
    assign pp1[2]   = a[2]  & b[1];
    assign pp2[2]   = a[2]  & b[2];
    assign pp3[2]   = a[2]  & b[3];
    assign pp4[2]   = a[2]  & b[4];
    assign pp5[2]   = a[2]  & b[5];
    assign pp6[2]   = a[2]  & b[6];
    assign pp7[2]   = a[2]  & b[7];
    assign pp8[2]   = a[2]  & b[8];
    assign pp9[2]   = a[2]  & b[9];
    assign pp10[2]  = a[2]  & b[10];
    assign pp11[2]  = a[2]  & b[11];
    assign pp12[2]  = a[2]  & b[12];
    assign pp13[2]  = a[2]  & b[13];
    assign pp14[2]  = a[2]  & b[14];
    assign pp15[2]  = a[2]  & b[15];
    assign pp16[2]  = a[2]  & b[16];
    assign pp17[2]  = a[2]  & b[17];
    assign pp18[2]  = a[2]  & b[18];
    assign pp19[2]  = a[2]  & b[19];
    assign pp20[2]  = a[2]  & b[20];
    assign pp21[2]  = a[2]  & b[21];
    assign pp22[2]  = a[2]  & b[22];
    assign pp23[2]  = a[2]  & b[23];
    assign pp24[2]  = a[2]  & b[24];
    assign pp25[2]  = a[2]  & b[25];
    assign pp26[2]  = a[2]  & b[26];
    assign pp27[2]  = a[2]  & b[27];
    assign pp28[2]  = a[2]  & b[28];
    assign pp29[2]  = a[2]  & b[29];
    assign pp30[2]  = a[2]  & b[30];
    assign pp31[2]  = a[2]  & b[31];

    assign pp0[3]   = a[3]  & b[0];
    assign pp1[3]   = a[3]  & b[1];
    assign pp2[3]   = a[3]  & b[2];
    assign pp3[3]   = a[3]  & b[3];
    assign pp4[3]   = a[3]  & b[4];
    assign pp5[3]   = a[3]  & b[5];
    assign pp6[3]   = a[3]  & b[6];
    assign pp7[3]   = a[3]  & b[7];
    assign pp8[3]   = a[3]  & b[8];
    assign pp9[3]   = a[3]  & b[9];
    assign pp10[3]  = a[3]  & b[10];
    assign pp11[3]  = a[3]  & b[11];
    assign pp12[3]  = a[3]  & b[12];
    assign pp13[3]  = a[3]  & b[13];
    assign pp14[3]  = a[3]  & b[14];
    assign pp15[3]  = a[3]  & b[15];
    assign pp16[3]  = a[3]  & b[16];
    assign pp17[3]  = a[3]  & b[17];
    assign pp18[3]  = a[3]  & b[18];
    assign pp19[3]  = a[3]  & b[19];
    assign pp20[3]  = a[3]  & b[20];
    assign pp21[3]  = a[3]  & b[21];
    assign pp22[3]  = a[3]  & b[22];
    assign pp23[3]  = a[3]  & b[23];
    assign pp24[3]  = a[3]  & b[24];
    assign pp25[3]  = a[3]  & b[25];
    assign pp26[3]  = a[3]  & b[26];
    assign pp27[3]  = a[3]  & b[27];
    assign pp28[3]  = a[3]  & b[28];
    assign pp29[3]  = a[3]  & b[29];
    assign pp30[3]  = a[3]  & b[30];
    assign pp31[3]  = a[3]  & b[31];

    assign pp0[4]   = a[4]  & b[0];
    assign pp1[4]   = a[4]  & b[1];
    assign pp2[4]   = a[4]  & b[2];
    assign pp3[4]   = a[4]  & b[3];
    assign pp4[4]   = a[4]  & b[4];
    assign pp5[4]   = a[4]  & b[5];
    assign pp6[4]   = a[4]  & b[6];
    assign pp7[4]   = a[4]  & b[7];
    assign pp8[4]   = a[4]  & b[8];
    assign pp9[4]   = a[4]  & b[9];
    assign pp10[4]  = a[4]  & b[10];
    assign pp11[4]  = a[4]  & b[11];
    assign pp12[4]  = a[4]  & b[12];
    assign pp13[4]  = a[4]  & b[13];
    assign pp14[4]  = a[4]  & b[14];
    assign pp15[4]  = a[4]  & b[15];
    assign pp16[4]  = a[4]  & b[16];
    assign pp17[4]  = a[4]  & b[17];
    assign pp18[4]  = a[4]  & b[18];
    assign pp19[4]  = a[4]  & b[19];
    assign pp20[4]  = a[4]  & b[20];
    assign pp21[4]  = a[4]  & b[21];
    assign pp22[4]  = a[4]  & b[22];
    assign pp23[4]  = a[4]  & b[23];
    assign pp24[4]  = a[4]  & b[24];
    assign pp25[4]  = a[4]  & b[25];
    assign pp26[4]  = a[4]  & b[26];
    assign pp27[4]  = a[4]  & b[27];
    assign pp28[4]  = a[4]  & b[28];
    assign pp29[4]  = a[4]  & b[29];
    assign pp30[4]  = a[4]  & b[30];
    assign pp31[4]  = a[4]  & b[31];

    assign pp0[5]   = a[5]  & b[0];
    assign pp1[5]   = a[5]  & b[1];
    assign pp2[5]   = a[5]  & b[2];
    assign pp3[5]   = a[5]  & b[3];
    assign pp4[5]   = a[5]  & b[4];
    assign pp5[5]   = a[5]  & b[5];
    assign pp6[5]   = a[5]  & b[6];
    assign pp7[5]   = a[5]  & b[7];
    assign pp8[5]   = a[5]  & b[8];
    assign pp9[5]   = a[5]  & b[9];
    assign pp10[5]  = a[5]  & b[10];
    assign pp11[5]  = a[5]  & b[11];
    assign pp12[5]  = a[5]  & b[12];
    assign pp13[5]  = a[5]  & b[13];
    assign pp14[5]  = a[5]  & b[14];
    assign pp15[5]  = a[5]  & b[15];
    assign pp16[5]  = a[5]  & b[16];
    assign pp17[5]  = a[5]  & b[17];
    assign pp18[5]  = a[5]  & b[18];
    assign pp19[5]  = a[5]  & b[19];
    assign pp20[5]  = a[5]  & b[20];
    assign pp21[5]  = a[5]  & b[21];
    assign pp22[5]  = a[5]  & b[22];
    assign pp23[5]  = a[5]  & b[23];
    assign pp24[5]  = a[5]  & b[24];
    assign pp25[5]  = a[5]  & b[25];
    assign pp26[5]  = a[5]  & b[26];
    assign pp27[5]  = a[5]  & b[27];
    assign pp28[5]  = a[5]  & b[28];
    assign pp29[5]  = a[5]  & b[29];
    assign pp30[5]  = a[5]  & b[30];
    assign pp31[5]  = a[5]  & b[31];

    assign pp0[6]   = a[6]  & b[0];
    assign pp1[6]   = a[6]  & b[1];
    assign pp2[6]   = a[6]  & b[2];
    assign pp3[6]   = a[6]  & b[3];
    assign pp4[6]   = a[6]  & b[4];
    assign pp5[6]   = a[6]  & b[5];
    assign pp6[6]   = a[6]  & b[6];
    assign pp7[6]   = a[6]  & b[7];
    assign pp8[6]   = a[6]  & b[8];
    assign pp9[6]   = a[6]  & b[9];
    assign pp10[6]  = a[6]  & b[10];
    assign pp11[6]  = a[6]  & b[11];
    assign pp12[6]  = a[6]  & b[12];
    assign pp13[6]  = a[6]  & b[13];
    assign pp14[6]  = a[6]  & b[14];
    assign pp15[6]  = a[6]  & b[15];
    assign pp16[6]  = a[6]  & b[16];
    assign pp17[6]  = a[6]  & b[17];
    assign pp18[6]  = a[6]  & b[18];
    assign pp19[6]  = a[6]  & b[19];
    assign pp20[6]  = a[6]  & b[20];
    assign pp21[6]  = a[6]  & b[21];
    assign pp22[6]  = a[6]  & b[22];
    assign pp23[6]  = a[6]  & b[23];
    assign pp24[6]  = a[6]  & b[24];
    assign pp25[6]  = a[6]  & b[25];
    assign pp26[6]  = a[6]  & b[26];
    assign pp27[6]  = a[6]  & b[27];
    assign pp28[6]  = a[6]  & b[28];
    assign pp29[6]  = a[6]  & b[29];
    assign pp30[6]  = a[6]  & b[30];
    assign pp31[6]  = a[6]  & b[31];

    assign pp0[7]   = a[7]  & b[0];
    assign pp1[7]   = a[7]  & b[1];
    assign pp2[7]   = a[7]  & b[2];
    assign pp3[7]   = a[7]  & b[3];
    assign pp4[7]   = a[7]  & b[4];
    assign pp5[7]   = a[7]  & b[5];
    assign pp6[7]   = a[7]  & b[6];
    assign pp7[7]   = a[7]  & b[7];
    assign pp8[7]   = a[7]  & b[8];
    assign pp9[7]   = a[7]  & b[9];
    assign pp10[7]  = a[7]  & b[10];
    assign pp11[7]  = a[7]  & b[11];
    assign pp12[7]  = a[7]  & b[12];
    assign pp13[7]  = a[7]  & b[13];
    assign pp14[7]  = a[7]  & b[14];
    assign pp15[7]  = a[7]  & b[15];
    assign pp16[7]  = a[7]  & b[16];
    assign pp17[7]  = a[7]  & b[17];
    assign pp18[7]  = a[7]  & b[18];
    assign pp19[7]  = a[7]  & b[19];
    assign pp20[7]  = a[7]  & b[20];
    assign pp21[7]  = a[7]  & b[21];
    assign pp22[7]  = a[7]  & b[22];
    assign pp23[7]  = a[7]  & b[23];
    assign pp24[7]  = a[7]  & b[24];
    assign pp25[7]  = a[7]  & b[25];
    assign pp26[7]  = a[7]  & b[26];
    assign pp27[7]  = a[7]  & b[27];
    assign pp28[7]  = a[7]  & b[28];
    assign pp29[7]  = a[7]  & b[29];
    assign pp30[7]  = a[7]  & b[30];
    assign pp31[7]  = a[7]  & b[31];

    assign pp0[8]   = a[8]  & b[0];
    assign pp1[8]   = a[8]  & b[1];
    assign pp2[8]   = a[8]  & b[2];
    assign pp3[8]   = a[8]  & b[3];
    assign pp4[8]   = a[8]  & b[4];
    assign pp5[8]   = a[8]  & b[5];
    assign pp6[8]   = a[8]  & b[6];
    assign pp7[8]   = a[8]  & b[7];
    assign pp8[8]   = a[8]  & b[8];
    assign pp9[8]   = a[8]  & b[9];
    assign pp10[8]  = a[8]  & b[10];
    assign pp11[8]  = a[8]  & b[11];
    assign pp12[8]  = a[8]  & b[12];
    assign pp13[8]  = a[8]  & b[13];
    assign pp14[8]  = a[8]  & b[14];
    assign pp15[8]  = a[8]  & b[15];
    assign pp16[8]  = a[8]  & b[16];
    assign pp17[8]  = a[8]  & b[17];
    assign pp18[8]  = a[8]  & b[18];
    assign pp19[8]  = a[8]  & b[19];
    assign pp20[8]  = a[8]  & b[20];
    assign pp21[8]  = a[8]  & b[21];
    assign pp22[8]  = a[8]  & b[22];
    assign pp23[8]  = a[8]  & b[23];
    assign pp24[8]  = a[8]  & b[24];
    assign pp25[8]  = a[8]  & b[25];
    assign pp26[8]  = a[8]  & b[26];
    assign pp27[8]  = a[8]  & b[27];
    assign pp28[8]  = a[8]  & b[28];
    assign pp29[8]  = a[8]  & b[29];
    assign pp30[8]  = a[8]  & b[30];
    assign pp31[8]  = a[8]  & b[31];

    assign pp0[9]   = a[9]  & b[0];
    assign pp1[9]   = a[9]  & b[1];
    assign pp2[9]   = a[9]  & b[2];
    assign pp3[9]   = a[9]  & b[3];
    assign pp4[9]   = a[9]  & b[4];
    assign pp5[9]   = a[9]  & b[5];
    assign pp6[9]   = a[9]  & b[6];
    assign pp7[9]   = a[9]  & b[7];
    assign pp8[9]   = a[9]  & b[8];
    assign pp9[9]   = a[9]  & b[9];
    assign pp10[9]  = a[9]  & b[10];
    assign pp11[9]  = a[9]  & b[11];
    assign pp12[9]  = a[9]  & b[12];
    assign pp13[9]  = a[9]  & b[13];
    assign pp14[9]  = a[9]  & b[14];
    assign pp15[9]  = a[9]  & b[15];
    assign pp16[9]  = a[9]  & b[16];
    assign pp17[9]  = a[9]  & b[17];
    assign pp18[9]  = a[9]  & b[18];
    assign pp19[9]  = a[9]  & b[19];
    assign pp20[9]  = a[9]  & b[20];
    assign pp21[9]  = a[9]  & b[21];
    assign pp22[9]  = a[9]  & b[22];
    assign pp23[9]  = a[9]  & b[23];
    assign pp24[9]  = a[9]  & b[24];
    assign pp25[9]  = a[9]  & b[25];
    assign pp26[9]  = a[9]  & b[26];
    assign pp27[9]  = a[9]  & b[27];
    assign pp28[9]  = a[9]  & b[28];
    assign pp29[9]  = a[9]  & b[29];
    assign pp30[9]  = a[9]  & b[30];
    assign pp31[9]  = a[9]  & b[31];

    assign pp0[10]   = a[10]  & b[0];
    assign pp1[10]   = a[10]  & b[1];
    assign pp2[10]   = a[10]  & b[2];
    assign pp3[10]   = a[10]  & b[3];
    assign pp4[10]   = a[10]  & b[4];
    assign pp5[10]   = a[10]  & b[5];
    assign pp6[10]   = a[10]  & b[6];
    assign pp7[10]   = a[10]  & b[7];
    assign pp8[10]   = a[10]  & b[8];
    assign pp9[10]   = a[10]  & b[9];
    assign pp10[10]  = a[10]  & b[10];
    assign pp11[10]  = a[10]  & b[11];
    assign pp12[10]  = a[10]  & b[12];
    assign pp13[10]  = a[10]  & b[13];
    assign pp14[10]  = a[10]  & b[14];
    assign pp15[10]  = a[10]  & b[15];
    assign pp16[10]  = a[10]  & b[16];
    assign pp17[10]  = a[10]  & b[17];
    assign pp18[10]  = a[10]  & b[18];
    assign pp19[10]  = a[10]  & b[19];
    assign pp20[10]  = a[10]  & b[20];
    assign pp21[10]  = a[10]  & b[21];
    assign pp22[10]  = a[10]  & b[22];
    assign pp23[10]  = a[10]  & b[23];
    assign pp24[10]  = a[10]  & b[24];
    assign pp25[10]  = a[10]  & b[25];
    assign pp26[10]  = a[10]  & b[26];
    assign pp27[10]  = a[10]  & b[27];
    assign pp28[10]  = a[10]  & b[28];
    assign pp29[10]  = a[10]  & b[29];
    assign pp30[10]  = a[10]  & b[30];
    assign pp31[10]  = a[10]  & b[31];

    assign pp0[11]   = a[11]  & b[0];
    assign pp1[11]   = a[11]  & b[1];
    assign pp2[11]   = a[11]  & b[2];
    assign pp3[11]   = a[11]  & b[3];
    assign pp4[11]   = a[11]  & b[4];
    assign pp5[11]   = a[11]  & b[5];
    assign pp6[11]   = a[11]  & b[6];
    assign pp7[11]   = a[11]  & b[7];
    assign pp8[11]   = a[11]  & b[8];
    assign pp9[11]   = a[11]  & b[9];
    assign pp10[11]  = a[11]  & b[10];
    assign pp11[11]  = a[11]  & b[11];
    assign pp12[11]  = a[11]  & b[12];
    assign pp13[11]  = a[11]  & b[13];
    assign pp14[11]  = a[11]  & b[14];
    assign pp15[11]  = a[11]  & b[15];
    assign pp16[11]  = a[11]  & b[16];
    assign pp17[11]  = a[11]  & b[17];
    assign pp18[11]  = a[11]  & b[18];
    assign pp19[11]  = a[11]  & b[19];
    assign pp20[11]  = a[11]  & b[20];
    assign pp21[11]  = a[11]  & b[21];
    assign pp22[11]  = a[11]  & b[22];
    assign pp23[11]  = a[11]  & b[23];
    assign pp24[11]  = a[11]  & b[24];
    assign pp25[11]  = a[11]  & b[25];
    assign pp26[11]  = a[11]  & b[26];
    assign pp27[11]  = a[11]  & b[27];
    assign pp28[11]  = a[11]  & b[28];
    assign pp29[11]  = a[11]  & b[29];
    assign pp30[11]  = a[11]  & b[30];
    assign pp31[11]  = a[11]  & b[31];

    assign pp0[12]   = a[12]  & b[0];
    assign pp1[12]   = a[12]  & b[1];
    assign pp2[12]   = a[12]  & b[2];
    assign pp3[12]   = a[12]  & b[3];
    assign pp4[12]   = a[12]  & b[4];
    assign pp5[12]   = a[12]  & b[5];
    assign pp6[12]   = a[12]  & b[6];
    assign pp7[12]   = a[12]  & b[7];
    assign pp8[12]   = a[12]  & b[8];
    assign pp9[12]   = a[12]  & b[9];
    assign pp10[12]  = a[12]  & b[10];
    assign pp11[12]  = a[12]  & b[11];
    assign pp12[12]  = a[12]  & b[12];
    assign pp13[12]  = a[12]  & b[13];
    assign pp14[12]  = a[12]  & b[14];
    assign pp15[12]  = a[12]  & b[15];
    assign pp16[12]  = a[12]  & b[16];
    assign pp17[12]  = a[12]  & b[17];
    assign pp18[12]  = a[12]  & b[18];
    assign pp19[12]  = a[12]  & b[19];
    assign pp20[12]  = a[12]  & b[20];
    assign pp21[12]  = a[12]  & b[21];
    assign pp22[12]  = a[12]  & b[22];
    assign pp23[12]  = a[12]  & b[23];
    assign pp24[12]  = a[12]  & b[24];
    assign pp25[12]  = a[12]  & b[25];
    assign pp26[12]  = a[12]  & b[26];
    assign pp27[12]  = a[12]  & b[27];
    assign pp28[12]  = a[12]  & b[28];
    assign pp29[12]  = a[12]  & b[29];
    assign pp30[12]  = a[12]  & b[30];
    assign pp31[12]  = a[12]  & b[31];

    assign pp0[13]   = a[13]  & b[0];
    assign pp1[13]   = a[13]  & b[1];
    assign pp2[13]   = a[13]  & b[2];
    assign pp3[13]   = a[13]  & b[3];
    assign pp4[13]   = a[13]  & b[4];
    assign pp5[13]   = a[13]  & b[5];
    assign pp6[13]   = a[13]  & b[6];
    assign pp7[13]   = a[13]  & b[7];
    assign pp8[13]   = a[13]  & b[8];
    assign pp9[13]   = a[13]  & b[9];
    assign pp10[13]  = a[13]  & b[10];
    assign pp11[13]  = a[13]  & b[11];
    assign pp12[13]  = a[13]  & b[12];
    assign pp13[13]  = a[13]  & b[13];
    assign pp14[13]  = a[13]  & b[14];
    assign pp15[13]  = a[13]  & b[15];
    assign pp16[13]  = a[13]  & b[16];
    assign pp17[13]  = a[13]  & b[17];
    assign pp18[13]  = a[13]  & b[18];
    assign pp19[13]  = a[13]  & b[19];
    assign pp20[13]  = a[13]  & b[20];
    assign pp21[13]  = a[13]  & b[21];
    assign pp22[13]  = a[13]  & b[22];
    assign pp23[13]  = a[13]  & b[23];
    assign pp24[13]  = a[13]  & b[24];
    assign pp25[13]  = a[13]  & b[25];
    assign pp26[13]  = a[13]  & b[26];
    assign pp27[13]  = a[13]  & b[27];
    assign pp28[13]  = a[13]  & b[28];
    assign pp29[13]  = a[13]  & b[29];
    assign pp30[13]  = a[13]  & b[30];
    assign pp31[13]  = a[13]  & b[31];

    assign pp0[14]   = a[14]  & b[0];
    assign pp1[14]   = a[14]  & b[1];
    assign pp2[14]   = a[14]  & b[2];
    assign pp3[14]   = a[14]  & b[3];
    assign pp4[14]   = a[14]  & b[4];
    assign pp5[14]   = a[14]  & b[5];
    assign pp6[14]   = a[14]  & b[6];
    assign pp7[14]   = a[14]  & b[7];
    assign pp8[14]   = a[14]  & b[8];
    assign pp9[14]   = a[14]  & b[9];
    assign pp10[14]  = a[14]  & b[10];
    assign pp11[14]  = a[14]  & b[11];
    assign pp12[14]  = a[14]  & b[12];
    assign pp13[14]  = a[14]  & b[13];
    assign pp14[14]  = a[14]  & b[14];
    assign pp15[14]  = a[14]  & b[15];
    assign pp16[14]  = a[14]  & b[16];
    assign pp17[14]  = a[14]  & b[17];
    assign pp18[14]  = a[14]  & b[18];
    assign pp19[14]  = a[14]  & b[19];
    assign pp20[14]  = a[14]  & b[20];
    assign pp21[14]  = a[14]  & b[21];
    assign pp22[14]  = a[14]  & b[22];
    assign pp23[14]  = a[14]  & b[23];
    assign pp24[14]  = a[14]  & b[24];
    assign pp25[14]  = a[14]  & b[25];
    assign pp26[14]  = a[14]  & b[26];
    assign pp27[14]  = a[14]  & b[27];
    assign pp28[14]  = a[14]  & b[28];
    assign pp29[14]  = a[14]  & b[29];
    assign pp30[14]  = a[14]  & b[30];
    assign pp31[14]  = a[14]  & b[31];

    assign pp0[15]   = a[15]  & b[0];
    assign pp1[15]   = a[15]  & b[1];
    assign pp2[15]   = a[15]  & b[2];
    assign pp3[15]   = a[15]  & b[3];
    assign pp4[15]   = a[15]  & b[4];
    assign pp5[15]   = a[15]  & b[5];
    assign pp6[15]   = a[15]  & b[6];
    assign pp7[15]   = a[15]  & b[7];
    assign pp8[15]   = a[15]  & b[8];
    assign pp9[15]   = a[15]  & b[9];
    assign pp10[15]  = a[15]  & b[10];
    assign pp11[15]  = a[15]  & b[11];
    assign pp12[15]  = a[15]  & b[12];
    assign pp13[15]  = a[15]  & b[13];
    assign pp14[15]  = a[15]  & b[14];
    assign pp15[15]  = a[15]  & b[15];
    assign pp16[15]  = a[15]  & b[16];
    assign pp17[15]  = a[15]  & b[17];
    assign pp18[15]  = a[15]  & b[18];
    assign pp19[15]  = a[15]  & b[19];
    assign pp20[15]  = a[15]  & b[20];
    assign pp21[15]  = a[15]  & b[21];
    assign pp22[15]  = a[15]  & b[22];
    assign pp23[15]  = a[15]  & b[23];
    assign pp24[15]  = a[15]  & b[24];
    assign pp25[15]  = a[15]  & b[25];
    assign pp26[15]  = a[15]  & b[26];
    assign pp27[15]  = a[15]  & b[27];
    assign pp28[15]  = a[15]  & b[28];
    assign pp29[15]  = a[15]  & b[29];
    assign pp30[15]  = a[15]  & b[30];
    assign pp31[15]  = a[15]  & b[31];

    assign pp0[16]   = a[16]  & b[0];
    assign pp1[16]   = a[16]  & b[1];
    assign pp2[16]   = a[16]  & b[2];
    assign pp3[16]   = a[16]  & b[3];
    assign pp4[16]   = a[16]  & b[4];
    assign pp5[16]   = a[16]  & b[5];
    assign pp6[16]   = a[16]  & b[6];
    assign pp7[16]   = a[16]  & b[7];
    assign pp8[16]   = a[16]  & b[8];
    assign pp9[16]   = a[16]  & b[9];
    assign pp10[16]  = a[16]  & b[10];
    assign pp11[16]  = a[16]  & b[11];
    assign pp12[16]  = a[16]  & b[12];
    assign pp13[16]  = a[16]  & b[13];
    assign pp14[16]  = a[16]  & b[14];
    assign pp15[16]  = a[16]  & b[15];
    assign pp16[16]  = a[16]  & b[16];
    assign pp17[16]  = a[16]  & b[17];
    assign pp18[16]  = a[16]  & b[18];
    assign pp19[16]  = a[16]  & b[19];
    assign pp20[16]  = a[16]  & b[20];
    assign pp21[16]  = a[16]  & b[21];
    assign pp22[16]  = a[16]  & b[22];
    assign pp23[16]  = a[16]  & b[23];
    assign pp24[16]  = a[16]  & b[24];
    assign pp25[16]  = a[16]  & b[25];
    assign pp26[16]  = a[16]  & b[26];
    assign pp27[16]  = a[16]  & b[27];
    assign pp28[16]  = a[16]  & b[28];
    assign pp29[16]  = a[16]  & b[29];
    assign pp30[16]  = a[16]  & b[30];
    assign pp31[16]  = a[16]  & b[31];

    assign pp0[17]   = a[17]  & b[0];
    assign pp1[17]   = a[17]  & b[1];
    assign pp2[17]   = a[17]  & b[2];
    assign pp3[17]   = a[17]  & b[3];
    assign pp4[17]   = a[17]  & b[4];
    assign pp5[17]   = a[17]  & b[5];
    assign pp6[17]   = a[17]  & b[6];
    assign pp7[17]   = a[17]  & b[7];
    assign pp8[17]   = a[17]  & b[8];
    assign pp9[17]   = a[17]  & b[9];
    assign pp10[17]  = a[17]  & b[10];
    assign pp11[17]  = a[17]  & b[11];
    assign pp12[17]  = a[17]  & b[12];
    assign pp13[17]  = a[17]  & b[13];
    assign pp14[17]  = a[17]  & b[14];
    assign pp15[17]  = a[17]  & b[15];
    assign pp16[17]  = a[17]  & b[16];
    assign pp17[17]  = a[17]  & b[17];
    assign pp18[17]  = a[17]  & b[18];
    assign pp19[17]  = a[17]  & b[19];
    assign pp20[17]  = a[17]  & b[20];
    assign pp21[17]  = a[17]  & b[21];
    assign pp22[17]  = a[17]  & b[22];
    assign pp23[17]  = a[17]  & b[23];
    assign pp24[17]  = a[17]  & b[24];
    assign pp25[17]  = a[17]  & b[25];
    assign pp26[17]  = a[17]  & b[26];
    assign pp27[17]  = a[17]  & b[27];
    assign pp28[17]  = a[17]  & b[28];
    assign pp29[17]  = a[17]  & b[29];
    assign pp30[17]  = a[17]  & b[30];
    assign pp31[17]  = a[17]  & b[31];

    assign pp0[18]   = a[18]  & b[0];
    assign pp1[18]   = a[18]  & b[1];
    assign pp2[18]   = a[18]  & b[2];
    assign pp3[18]   = a[18]  & b[3];
    assign pp4[18]   = a[18]  & b[4];
    assign pp5[18]   = a[18]  & b[5];
    assign pp6[18]   = a[18]  & b[6];
    assign pp7[18]   = a[18]  & b[7];
    assign pp8[18]   = a[18]  & b[8];
    assign pp9[18]   = a[18]  & b[9];
    assign pp10[18]  = a[18]  & b[10];
    assign pp11[18]  = a[18]  & b[11];
    assign pp12[18]  = a[18]  & b[12];
    assign pp13[18]  = a[18]  & b[13];
    assign pp14[18]  = a[18]  & b[14];
    assign pp15[18]  = a[18]  & b[15];
    assign pp16[18]  = a[18]  & b[16];
    assign pp17[18]  = a[18]  & b[17];
    assign pp18[18]  = a[18]  & b[18];
    assign pp19[18]  = a[18]  & b[19];
    assign pp20[18]  = a[18]  & b[20];
    assign pp21[18]  = a[18]  & b[21];
    assign pp22[18]  = a[18]  & b[22];
    assign pp23[18]  = a[18]  & b[23];
    assign pp24[18]  = a[18]  & b[24];
    assign pp25[18]  = a[18]  & b[25];
    assign pp26[18]  = a[18]  & b[26];
    assign pp27[18]  = a[18]  & b[27];
    assign pp28[18]  = a[18]  & b[28];
    assign pp29[18]  = a[18]  & b[29];
    assign pp30[18]  = a[18]  & b[30];
    assign pp31[18]  = a[18]  & b[31];

    assign pp0[19]   = a[19]  & b[0];
    assign pp1[19]   = a[19]  & b[1];
    assign pp2[19]   = a[19]  & b[2];
    assign pp3[19]   = a[19]  & b[3];
    assign pp4[19]   = a[19]  & b[4];
    assign pp5[19]   = a[19]  & b[5];
    assign pp6[19]   = a[19]  & b[6];
    assign pp7[19]   = a[19]  & b[7];
    assign pp8[19]   = a[19]  & b[8];
    assign pp9[19]   = a[19]  & b[9];
    assign pp10[19]  = a[19]  & b[10];
    assign pp11[19]  = a[19]  & b[11];
    assign pp12[19]  = a[19]  & b[12];
    assign pp13[19]  = a[19]  & b[13];
    assign pp14[19]  = a[19]  & b[14];
    assign pp15[19]  = a[19]  & b[15];
    assign pp16[19]  = a[19]  & b[16];
    assign pp17[19]  = a[19]  & b[17];
    assign pp18[19]  = a[19]  & b[18];
    assign pp19[19]  = a[19]  & b[19];
    assign pp20[19]  = a[19]  & b[20];
    assign pp21[19]  = a[19]  & b[21];
    assign pp22[19]  = a[19]  & b[22];
    assign pp23[19]  = a[19]  & b[23];
    assign pp24[19]  = a[19]  & b[24];
    assign pp25[19]  = a[19]  & b[25];
    assign pp26[19]  = a[19]  & b[26];
    assign pp27[19]  = a[19]  & b[27];
    assign pp28[19]  = a[19]  & b[28];
    assign pp29[19]  = a[19]  & b[29];
    assign pp30[19]  = a[19]  & b[30];
    assign pp31[19]  = a[19]  & b[31];

    assign pp0[20]   = a[20]  & b[0];
    assign pp1[20]   = a[20]  & b[1];
    assign pp2[20]   = a[20]  & b[2];
    assign pp3[20]   = a[20]  & b[3];
    assign pp4[20]   = a[20]  & b[4];
    assign pp5[20]   = a[20]  & b[5];
    assign pp6[20]   = a[20]  & b[6];
    assign pp7[20]   = a[20]  & b[7];
    assign pp8[20]   = a[20]  & b[8];
    assign pp9[20]   = a[20]  & b[9];
    assign pp10[20]  = a[20]  & b[10];
    assign pp11[20]  = a[20]  & b[11];
    assign pp12[20]  = a[20]  & b[12];
    assign pp13[20]  = a[20]  & b[13];
    assign pp14[20]  = a[20]  & b[14];
    assign pp15[20]  = a[20]  & b[15];
    assign pp16[20]  = a[20]  & b[16];
    assign pp17[20]  = a[20]  & b[17];
    assign pp18[20]  = a[20]  & b[18];
    assign pp19[20]  = a[20]  & b[19];
    assign pp20[20]  = a[20]  & b[20];
    assign pp21[20]  = a[20]  & b[21];
    assign pp22[20]  = a[20]  & b[22];
    assign pp23[20]  = a[20]  & b[23];
    assign pp24[20]  = a[20]  & b[24];
    assign pp25[20]  = a[20]  & b[25];
    assign pp26[20]  = a[20]  & b[26];
    assign pp27[20]  = a[20]  & b[27];
    assign pp28[20]  = a[20]  & b[28];
    assign pp29[20]  = a[20]  & b[29];
    assign pp30[20]  = a[20]  & b[30];
    assign pp31[20]  = a[20]  & b[31];

    assign pp0[21]   = a[21]  & b[0];
    assign pp1[21]   = a[21]  & b[1];
    assign pp2[21]   = a[21]  & b[2];
    assign pp3[21]   = a[21]  & b[3];
    assign pp4[21]   = a[21]  & b[4];
    assign pp5[21]   = a[21]  & b[5];
    assign pp6[21]   = a[21]  & b[6];
    assign pp7[21]   = a[21]  & b[7];
    assign pp8[21]   = a[21]  & b[8];
    assign pp9[21]   = a[21]  & b[9];
    assign pp10[21]  = a[21]  & b[10];
    assign pp11[21]  = a[21]  & b[11];
    assign pp12[21]  = a[21]  & b[12];
    assign pp13[21]  = a[21]  & b[13];
    assign pp14[21]  = a[21]  & b[14];
    assign pp15[21]  = a[21]  & b[15];
    assign pp16[21]  = a[21]  & b[16];
    assign pp17[21]  = a[21]  & b[17];
    assign pp18[21]  = a[21]  & b[18];
    assign pp19[21]  = a[21]  & b[19];
    assign pp20[21]  = a[21]  & b[20];
    assign pp21[21]  = a[21]  & b[21];
    assign pp22[21]  = a[21]  & b[22];
    assign pp23[21]  = a[21]  & b[23];
    assign pp24[21]  = a[21]  & b[24];
    assign pp25[21]  = a[21]  & b[25];
    assign pp26[21]  = a[21]  & b[26];
    assign pp27[21]  = a[21]  & b[27];
    assign pp28[21]  = a[21]  & b[28];
    assign pp29[21]  = a[21]  & b[29];
    assign pp30[21]  = a[21]  & b[30];
    assign pp31[21]  = a[21]  & b[31];
      
    assign pp0[22]   = a[22]  & b[0];
    assign pp1[22]   = a[22]  & b[1];
    assign pp2[22]   = a[22]  & b[2];
    assign pp3[22]   = a[22]  & b[3];
    assign pp4[22]   = a[22]  & b[4];
    assign pp5[22]   = a[22]  & b[5];
    assign pp6[22]   = a[22]  & b[6];
    assign pp7[22]   = a[22]  & b[7];
    assign pp8[22]   = a[22]  & b[8];
    assign pp9[22]   = a[22]  & b[9];
    assign pp10[22]  = a[22]  & b[10];
    assign pp11[22]  = a[22]  & b[11];
    assign pp12[22]  = a[22]  & b[12];
    assign pp13[22]  = a[22]  & b[13];
    assign pp14[22]  = a[22]  & b[14];
    assign pp15[22]  = a[22]  & b[15];
    assign pp16[22]  = a[22]  & b[16];
    assign pp17[22]  = a[22]  & b[17];
    assign pp18[22]  = a[22]  & b[18];
    assign pp19[22]  = a[22]  & b[19];
    assign pp20[22]  = a[22]  & b[20];
    assign pp21[22]  = a[22]  & b[21];
    assign pp22[22]  = a[22]  & b[22];
    assign pp23[22]  = a[22]  & b[23];
    assign pp24[22]  = a[22]  & b[24];
    assign pp25[22]  = a[22]  & b[25];
    assign pp26[22]  = a[22]  & b[26];
    assign pp27[22]  = a[22]  & b[27];
    assign pp28[22]  = a[22]  & b[28];
    assign pp29[22]  = a[22]  & b[29];
    assign pp30[22]  = a[22]  & b[30];
    assign pp31[22]  = a[22]  & b[31];

    assign pp0[23]   = a[23]  & b[0];
    assign pp1[23]   = a[23]  & b[1];
    assign pp2[23]   = a[23]  & b[2];
    assign pp3[23]   = a[23]  & b[3];
    assign pp4[23]   = a[23]  & b[4];
    assign pp5[23]   = a[23]  & b[5];
    assign pp6[23]   = a[23]  & b[6];
    assign pp7[23]   = a[23]  & b[7];
    assign pp8[23]   = a[23]  & b[8];
    assign pp9[23]   = a[23]  & b[9];
    assign pp10[23]  = a[23]  & b[10];
    assign pp11[23]  = a[23]  & b[11];
    assign pp12[23]  = a[23]  & b[12];
    assign pp13[23]  = a[23]  & b[13];
    assign pp14[23]  = a[23]  & b[14];
    assign pp15[23]  = a[23]  & b[15];
    assign pp16[23]  = a[23]  & b[16];
    assign pp17[23]  = a[23]  & b[17];
    assign pp18[23]  = a[23]  & b[18];
    assign pp19[23]  = a[23]  & b[19];
    assign pp20[23]  = a[23]  & b[20];
    assign pp21[23]  = a[23]  & b[21];
    assign pp22[23]  = a[23]  & b[22];
    assign pp23[23]  = a[23]  & b[23];
    assign pp24[23]  = a[23]  & b[24];
    assign pp25[23]  = a[23]  & b[25];
    assign pp26[23]  = a[23]  & b[26];
    assign pp27[23]  = a[23]  & b[27];
    assign pp28[23]  = a[23]  & b[28];
    assign pp29[23]  = a[23]  & b[29];
    assign pp30[23]  = a[23]  & b[30];
    assign pp31[23]  = a[23]  & b[31];

    assign pp0[24]   = a[24]  & b[0];
    assign pp1[24]   = a[24]  & b[1];
    assign pp2[24]   = a[24]  & b[2];
    assign pp3[24]   = a[24]  & b[3];
    assign pp4[24]   = a[24]  & b[4];
    assign pp5[24]   = a[24]  & b[5];
    assign pp6[24]   = a[24]  & b[6];
    assign pp7[24]   = a[24]  & b[7];
    assign pp8[24]   = a[24]  & b[8];
    assign pp9[24]   = a[24]  & b[9];
    assign pp10[24]  = a[24]  & b[10];
    assign pp11[24]  = a[24]  & b[11];
    assign pp12[24]  = a[24]  & b[12];
    assign pp13[24]  = a[24]  & b[13];
    assign pp14[24]  = a[24]  & b[14];
    assign pp15[24]  = a[24]  & b[15];
    assign pp16[24]  = a[24]  & b[16];
    assign pp17[24]  = a[24]  & b[17];
    assign pp18[24]  = a[24]  & b[18];
    assign pp19[24]  = a[24]  & b[19];
    assign pp20[24]  = a[24]  & b[20];
    assign pp21[24]  = a[24]  & b[21];
    assign pp22[24]  = a[24]  & b[22];
    assign pp23[24]  = a[24]  & b[23];
    assign pp24[24]  = a[24]  & b[24];
    assign pp25[24]  = a[24]  & b[25];
    assign pp26[24]  = a[24]  & b[26];
    assign pp27[24]  = a[24]  & b[27];
    assign pp28[24]  = a[24]  & b[28];
    assign pp29[24]  = a[24]  & b[29];
    assign pp30[24]  = a[24]  & b[30];
    assign pp31[24]  = a[24]  & b[31];

    assign pp0[25]   = a[25]  & b[0];
    assign pp1[25]   = a[25]  & b[1];
    assign pp2[25]   = a[25]  & b[2];
    assign pp3[25]   = a[25]  & b[3];
    assign pp4[25]   = a[25]  & b[4];
    assign pp5[25]   = a[25]  & b[5];
    assign pp6[25]   = a[25]  & b[6];
    assign pp7[25]   = a[25]  & b[7];
    assign pp8[25]   = a[25]  & b[8];
    assign pp9[25]   = a[25]  & b[9];
    assign pp10[25]  = a[25]  & b[10];
    assign pp11[25]  = a[25]  & b[11];
    assign pp12[25]  = a[25]  & b[12];
    assign pp13[25]  = a[25]  & b[13];
    assign pp14[25]  = a[25]  & b[14];
    assign pp15[25]  = a[25]  & b[15];
    assign pp16[25]  = a[25]  & b[16];
    assign pp17[25]  = a[25]  & b[17];
    assign pp18[25]  = a[25]  & b[18];
    assign pp19[25]  = a[25]  & b[19];
    assign pp20[25]  = a[25]  & b[20];
    assign pp21[25]  = a[25]  & b[21];
    assign pp22[25]  = a[25]  & b[22];
    assign pp23[25]  = a[25]  & b[23];
    assign pp24[25]  = a[25]  & b[24];
    assign pp25[25]  = a[25]  & b[25];
    assign pp26[25]  = a[25]  & b[26];
    assign pp27[25]  = a[25]  & b[27];
    assign pp28[25]  = a[25]  & b[28];
    assign pp29[25]  = a[25]  & b[29];
    assign pp30[25]  = a[25]  & b[30];
    assign pp31[25]  = a[25]  & b[31];

    assign pp0[26]   = a[26]  & b[0];
    assign pp1[26]   = a[26]  & b[1];
    assign pp2[26]   = a[26]  & b[2];
    assign pp3[26]   = a[26]  & b[3];
    assign pp4[26]   = a[26]  & b[4];
    assign pp5[26]   = a[26]  & b[5];
    assign pp6[26]   = a[26]  & b[6];
    assign pp7[26]   = a[26]  & b[7];
    assign pp8[26]   = a[26]  & b[8];
    assign pp9[26]   = a[26]  & b[9];
    assign pp10[26]  = a[26]  & b[10];
    assign pp11[26]  = a[26]  & b[11];
    assign pp12[26]  = a[26]  & b[12];
    assign pp13[26]  = a[26]  & b[13];
    assign pp14[26]  = a[26]  & b[14];
    assign pp15[26]  = a[26]  & b[15];
    assign pp16[26]  = a[26]  & b[16];
    assign pp17[26]  = a[26]  & b[17];
    assign pp18[26]  = a[26]  & b[18];
    assign pp19[26]  = a[26]  & b[19];
    assign pp20[26]  = a[26]  & b[20];
    assign pp21[26]  = a[26]  & b[21];
    assign pp22[26]  = a[26]  & b[22];
    assign pp23[26]  = a[26]  & b[23];
    assign pp24[26]  = a[26]  & b[24];
    assign pp25[26]  = a[26]  & b[25];
    assign pp26[26]  = a[26]  & b[26];
    assign pp27[26]  = a[26]  & b[27];
    assign pp28[26]  = a[26]  & b[28];
    assign pp29[26]  = a[26]  & b[29];
    assign pp30[26]  = a[26]  & b[30];
    assign pp31[26]  = a[26]  & b[31];

    assign pp0[27]   = a[27]  & b[0];
    assign pp1[27]   = a[27]  & b[1];
    assign pp2[27]   = a[27]  & b[2];
    assign pp3[27]   = a[27]  & b[3];
    assign pp4[27]   = a[27]  & b[4];
    assign pp5[27]   = a[27]  & b[5];
    assign pp6[27]   = a[27]  & b[6];
    assign pp7[27]   = a[27]  & b[7];
    assign pp8[27]   = a[27]  & b[8];
    assign pp9[27]   = a[27]  & b[9];
    assign pp10[27]  = a[27]  & b[10];
    assign pp11[27]  = a[27]  & b[11];
    assign pp12[27]  = a[27]  & b[12];
    assign pp13[27]  = a[27]  & b[13];
    assign pp14[27]  = a[27]  & b[14];
    assign pp15[27]  = a[27]  & b[15];
    assign pp16[27]  = a[27]  & b[16];
    assign pp17[27]  = a[27]  & b[17];
    assign pp18[27]  = a[27]  & b[18];
    assign pp19[27]  = a[27]  & b[19];
    assign pp20[27]  = a[27]  & b[20];
    assign pp21[27]  = a[27]  & b[21];
    assign pp22[27]  = a[27]  & b[22];
    assign pp23[27]  = a[27]  & b[23];
    assign pp24[27]  = a[27]  & b[24];
    assign pp25[27]  = a[27]  & b[25];
    assign pp26[27]  = a[27]  & b[26];
    assign pp27[27]  = a[27]  & b[27];
    assign pp28[27]  = a[27]  & b[28];
    assign pp29[27]  = a[27]  & b[29];
    assign pp30[27]  = a[27]  & b[30];
    assign pp31[27]  = a[27]  & b[31];

    assign pp0[28]   = a[28]  & b[0];
    assign pp1[28]   = a[28]  & b[1];
    assign pp2[28]   = a[28]  & b[2];
    assign pp3[28]   = a[28]  & b[3];
    assign pp4[28]   = a[28]  & b[4];
    assign pp5[28]   = a[28]  & b[5];
    assign pp6[28]   = a[28]  & b[6];
    assign pp7[28]   = a[28]  & b[7];
    assign pp8[28]   = a[28]  & b[8];
    assign pp9[28]   = a[28]  & b[9];
    assign pp10[28]  = a[28]  & b[10];
    assign pp11[28]  = a[28]  & b[11];
    assign pp12[28]  = a[28]  & b[12];
    assign pp13[28]  = a[28]  & b[13];
    assign pp14[28]  = a[28]  & b[14];
    assign pp15[28]  = a[28]  & b[15];
    assign pp16[28]  = a[28]  & b[16];
    assign pp17[28]  = a[28]  & b[17];
    assign pp18[28]  = a[28]  & b[18];
    assign pp19[28]  = a[28]  & b[19];
    assign pp20[28]  = a[28]  & b[20];
    assign pp21[28]  = a[28]  & b[21];
    assign pp22[28]  = a[28]  & b[22];
    assign pp23[28]  = a[28]  & b[23];
    assign pp24[28]  = a[28]  & b[24];
    assign pp25[28]  = a[28]  & b[25];
    assign pp26[28]  = a[28]  & b[26];
    assign pp27[28]  = a[28]  & b[27];
    assign pp28[28]  = a[28]  & b[28];
    assign pp29[28]  = a[28]  & b[29];
    assign pp30[28]  = a[28]  & b[30];
    assign pp31[28]  = a[28]  & b[31];

    assign pp0[29]   = a[29]  & b[0];
    assign pp1[29]   = a[29]  & b[1];
    assign pp2[29]   = a[29]  & b[2];
    assign pp3[29]   = a[29]  & b[3];
    assign pp4[29]   = a[29]  & b[4];
    assign pp5[29]   = a[29]  & b[5];
    assign pp6[29]   = a[29]  & b[6];
    assign pp7[29]   = a[29]  & b[7];
    assign pp8[29]   = a[29]  & b[8];
    assign pp9[29]   = a[29]  & b[9];
    assign pp10[29]  = a[29]  & b[10];
    assign pp11[29]  = a[29]  & b[11];
    assign pp12[29]  = a[29]  & b[12];
    assign pp13[29]  = a[29]  & b[13];
    assign pp14[29]  = a[29]  & b[14];
    assign pp15[29]  = a[29]  & b[15];
    assign pp16[29]  = a[29]  & b[16];
    assign pp17[29]  = a[29]  & b[17];
    assign pp18[29]  = a[29]  & b[18];
    assign pp19[29]  = a[29]  & b[19];
    assign pp20[29]  = a[29]  & b[20];
    assign pp21[29]  = a[29]  & b[21];
    assign pp22[29]  = a[29]  & b[22];
    assign pp23[29]  = a[29]  & b[23];
    assign pp24[29]  = a[29]  & b[24];
    assign pp25[29]  = a[29]  & b[25];
    assign pp26[29]  = a[29]  & b[26];
    assign pp27[29]  = a[29]  & b[27];
    assign pp28[29]  = a[29]  & b[28];
    assign pp29[29]  = a[29]  & b[29];
    assign pp30[29]  = a[29]  & b[30];
    assign pp31[29]  = a[29]  & b[31];

    assign pp0[30]   = a[30]  & b[0];
    assign pp1[30]   = a[30]  & b[1];
    assign pp2[30]   = a[30]  & b[2];
    assign pp3[30]   = a[30]  & b[3];
    assign pp4[30]   = a[30]  & b[4];
    assign pp5[30]   = a[30]  & b[5];
    assign pp6[30]   = a[30]  & b[6];
    assign pp7[30]   = a[30]  & b[7];
    assign pp8[30]   = a[30]  & b[8];
    assign pp9[30]   = a[30]  & b[9];
    assign pp10[30]  = a[30]  & b[10];
    assign pp11[30]  = a[30]  & b[11];
    assign pp12[30]  = a[30]  & b[12];
    assign pp13[30]  = a[30]  & b[13];
    assign pp14[30]  = a[30]  & b[14];
    assign pp15[30]  = a[30]  & b[15];
    assign pp16[30]  = a[30]  & b[16];
    assign pp17[30]  = a[30]  & b[17];
    assign pp18[30]  = a[30]  & b[18];
    assign pp19[30]  = a[30]  & b[19];
    assign pp20[30]  = a[30]  & b[20];
    assign pp21[30]  = a[30]  & b[21];
    assign pp22[30]  = a[30]  & b[22];
    assign pp23[30]  = a[30]  & b[23];
    assign pp24[30]  = a[30]  & b[24];
    assign pp25[30]  = a[30]  & b[25];
    assign pp26[30]  = a[30]  & b[26];
    assign pp27[30]  = a[30]  & b[27];
    assign pp28[30]  = a[30]  & b[28];
    assign pp29[30]  = a[30]  & b[29];
    assign pp30[30]  = a[30]  & b[30];
    assign pp31[30]  = a[30]  & b[31];

    assign pp0[31]   = a[31]  & b[0];
    assign pp1[31]   = a[31]  & b[1];
    assign pp2[31]   = a[31]  & b[2];
    assign pp3[31]   = a[31]  & b[3];
    assign pp4[31]   = a[31]  & b[4];
    assign pp5[31]   = a[31]  & b[5];
    assign pp6[31]   = a[31]  & b[6];
    assign pp7[31]   = a[31]  & b[7];
    assign pp8[31]   = a[31]  & b[8];
    assign pp9[31]   = a[31]  & b[9];
    assign pp10[31]  = a[31]  & b[10];
    assign pp11[31]  = a[31]  & b[11];
    assign pp12[31]  = a[31]  & b[12];
    assign pp13[31]  = a[31]  & b[13];
    assign pp14[31]  = a[31]  & b[14];
    assign pp15[31]  = a[31]  & b[15];
    assign pp16[31]  = a[31]  & b[16];
    assign pp17[31]  = a[31]  & b[17];
    assign pp18[31]  = a[31]  & b[18];
    assign pp19[31]  = a[31]  & b[19];
    assign pp20[31]  = a[31]  & b[20];
    assign pp21[31]  = a[31]  & b[21];
    assign pp22[31]  = a[31]  & b[22];
    assign pp23[31]  = a[31]  & b[23];
    assign pp24[31]  = a[31]  & b[24];
    assign pp25[31]  = a[31]  & b[25];
    assign pp26[31]  = a[31]  & b[26];
    assign pp27[31]  = a[31]  & b[27];
    assign pp28[31]  = a[31]  & b[28];
    assign pp29[31]  = a[31]  & b[29];
    assign pp30[31]  = a[31]  & b[30];
    assign pp31[31]  = a[31]  & b[31];

    // Template for Find & Replace
    // assign pp0[%]   = a[%]  & b[0];
    // assign pp1[%]   = a[%]  & b[1];
    // assign pp2[%]   = a[%]  & b[2];
    // assign pp3[%]   = a[%]  & b[3];
    // assign pp4[%]   = a[%]  & b[4];
    // assign pp5[%]   = a[%]  & b[5];
    // assign pp6[%]   = a[%]  & b[6];
    // assign pp7[%]   = a[%]  & b[7];
    // assign pp8[%]   = a[%]  & b[8];
    // assign pp9[%]   = a[%]  & b[9];
    // assign pp10[%]  = a[%]  & b[10];
    // assign pp11[%]  = a[%]  & b[11];
    // assign pp12[%]  = a[%]  & b[12];
    // assign pp13[%]  = a[%]  & b[13];
    // assign pp14[%]  = a[%]  & b[14];
    // assign pp15[%]  = a[%]  & b[15];
    // assign pp16[%]  = a[%]  & b[16];
    // assign pp17[%]  = a[%]  & b[17];
    // assign pp18[%]  = a[%]  & b[18];
    // assign pp19[%]  = a[%]  & b[19];
    // assign pp20[%]  = a[%]  & b[20];
    // assign pp21[%]  = a[%]  & b[21];
    // assign pp22[%]  = a[%]  & b[22];
    // assign pp23[%]  = a[%]  & b[23];
    // assign pp24[%]  = a[%]  & b[24];
    // assign pp25[%]  = a[%]  & b[25];
    // assign pp26[%]  = a[%]  & b[26];
    // assign pp27[%]  = a[%]  & b[27];
    // assign pp28[%]  = a[%]  & b[28];
    // assign pp29[%]  = a[%]  & b[29];
    // assign pp30[%]  = a[%]  & b[30];
    // assign pp31[%]  = a[%]  & b[31];
endmodule 
