// Compiler Directives

// Used for extra debug outputs for the LED display, turn on for FPGA prototyping, off for simulation
`define VALIDATION 1

// Used for pipeline testebenching, turn on to clock 5 times, off to clock once
`define PIPELINE 1